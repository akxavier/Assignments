module xor_gate
(output out,
input a, b);

xor g1 (out, a, b);

endmodule
module and_gate 
(output out,
input a, b);

and g1 (out, a, b);

endmodule
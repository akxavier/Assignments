module not_gate
(output x,
input y);

not g1 (x, y);

endmodule 
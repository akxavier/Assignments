module mult_signed(out, X, Y);

output [7:0] out;
input [3:0] X, Y;

assign out[0] = X[0] * Y[0],
	out [1] = (X[1] * Y[0]) + (X[0] * Y[1]),
	out [2] = (X[2] * Y[0]) + (X[1] * Y[1]) + (X[0] * Y[2]),
	out [3] = (X[3] * Y[0]) + (X[2] * Y[1]) + (X[1] * Y[2]) - (X[0] * Y[3]),
	out [4] = (X[3] * Y[0]) + (X[3] * Y[1]) + (X[2] * Y[2]) - (X[1] * Y[3]),
	out [5] = (X[3] * Y[0]) + (X[3] * Y[1]) + (X[3] * Y[2]) - (X[2] * Y[3]),
	out [6] = (X[3] * Y[0]) + (X[3] * Y[1]) + (X[3] * Y[2]) - (X[3] * Y[3]),
	out [7] = (X[3] * Y[0]) + (X[3] * Y[1]) + (X[3] * Y[2]) - (X[3] * Y[3]);
	
endmodule
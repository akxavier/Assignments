module array_of_16_inverters_gate 
(output [15:0] out,
input [15:0] in);

not g[15:0] (out, in);

endmodule
module array_of_16_and_gate
(output [15:0] out,
input [15:0] a, b);

and g[15:0] (out, a, b);

endmodule
module not_dataflow (out, in);

output out;
input in;

assign out = ~in;

endmodule
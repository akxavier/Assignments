module ripple_carry_dataflow32_tb;

wire [31:0] s;
wire cout;
reg [31:0] a, b;

ripple_carry_dataflow32 a1 (.s(s), .cout(cout), .a(a), .b(b));

initial 
begin
	a = 32'b00000000100000000000100000000000; b = 32'b00000000000000100000000000000000;
	#5 a = 32'b00000000100000000000000000000000; b = 32'b00000000000100000000000000000000;
	#5 a = 32'b00000000000000000000100000001000; b = 32'b00000000000010000000000000000000;
	#5 a = 32'b00000010000000000000100000000000; b = 32'b00000000000000000000000010000000;
	#5 a = 32'b00000000000000000100000000000000; b = 32'b00010000000000000000000000000000;
	#5 a = 32'b00000000001000000000000000100000; b = 32'b00000000000000000000001000000000;
	#5 a = 32'b00000000000011100000000000000000; b = 32'b00000000000000100000000000000000;
	#5 a = 32'b00000000000000000000100000000000; b = 32'b00100000000000000000000001000000;
	#5 a = 32'b00000001000000000000000000000000; b = 32'b00000000001000000011100000000000;
end

initial
$monitor ($time, "a = %b, b = %b, cout = %b, s = %b", a, b, cout, s);

endmodule
module xnor_gate
(output out,
input a, b);

xnor g1 (out, a, b);

endmodule 
module ripple_carry_dataflow32 (s, cout, a, b);

output [31:0] s;
output cout;
input [31:0] a, b;

wire [30:0] c;

fa_dataflow g0 (.s(s[0]), .cout(c[0]), .a(a[0]), .b(b[0]), .c(1'b0));
fa_dataflow g1 (.s(s[1]), .cout(c[1]), .a(a[1]), .b(b[1]), .c(c[0]));
fa_dataflow g2 (.s(s[2]), .cout(c[2]), .a(a[2]), .b(b[2]), .c(c[1]));
fa_dataflow g3 (.s(s[3]), .cout(c[3]), .a(a[3]), .b(b[3]), .c(c[2]));
fa_dataflow g4 (.s(s[4]), .cout(c[4]), .a(a[4]), .b(b[4]), .c(c[3]));
fa_dataflow g5 (.s(s[5]), .cout(c[5]), .a(a[5]), .b(b[5]), .c(c[4]));
fa_dataflow g6 (.s(s[6]), .cout(c[6]), .a(a[6]), .b(b[6]), .c(c[5]));
fa_dataflow g7 (.s(s[7]), .cout(c[7]), .a(a[7]), .b(b[7]), .c(c[6]));
fa_dataflow g8 (.s(s[8]), .cout(c[8]), .a(a[8]), .b(b[8]), .c(c[7]));
fa_dataflow g9 (.s(s[9]), .cout(c[9]), .a(a[9]), .b(b[9]), .c(c[8]));
fa_dataflow g10 (.s(s[10]), .cout(c[10]), .a(a[10]), .b(b[10]), .c(c[9]));
fa_dataflow g11 (.s(s[11]), .cout(c[11]), .a(a[11]), .b(b[11]), .c(c[10]));
fa_dataflow g12 (.s(s[12]), .cout(c[12]), .a(a[12]), .b(b[12]), .c(c[11]));
fa_dataflow g13 (.s(s[13]), .cout(c[13]), .a(a[13]), .b(b[13]), .c(c[12]));
fa_dataflow g14 (.s(s[14]), .cout(c[14]), .a(a[14]), .b(b[14]), .c(c[13]));
fa_dataflow g15 (.s(s[15]), .cout(c[15]), .a(a[15]), .b(b[15]), .c(c[14]));
fa_dataflow g16 (.s(s[16]), .cout(c[16]), .a(a[16]), .b(b[16]), .c(c[15]));
fa_dataflow g17 (.s(s[17]), .cout(c[17]), .a(a[17]), .b(b[17]), .c(c[16]));
fa_dataflow g18 (.s(s[18]), .cout(c[18]), .a(a[18]), .b(b[18]), .c(c[17]));
fa_dataflow g19 (.s(s[19]), .cout(c[19]), .a(a[19]), .b(b[19]), .c(c[18]));
fa_dataflow g20 (.s(s[20]), .cout(c[20]), .a(a[20]), .b(b[20]), .c(c[19]));
fa_dataflow g21 (.s(s[21]), .cout(c[21]), .a(a[21]), .b(b[21]), .c(c[20]));
fa_dataflow g22 (.s(s[22]), .cout(c[22]), .a(a[22]), .b(b[22]), .c(c[21]));
fa_dataflow g23 (.s(s[23]), .cout(c[23]), .a(a[23]), .b(b[23]), .c(c[22]));
fa_dataflow g24 (.s(s[24]), .cout(c[24]), .a(a[24]), .b(b[24]), .c(c[23]));
fa_dataflow g25 (.s(s[25]), .cout(c[25]), .a(a[25]), .b(b[25]), .c(c[24]));
fa_dataflow g26 (.s(s[26]), .cout(c[26]), .a(a[26]), .b(b[26]), .c(c[25]));
fa_dataflow g27 (.s(s[27]), .cout(c[27]), .a(a[27]), .b(b[27]), .c(c[26]));
fa_dataflow g28 (.s(s[28]), .cout(c[28]), .a(a[28]), .b(b[28]), .c(c[27]));
fa_dataflow g29 (.s(s[29]), .cout(c[29]), .a(a[29]), .b(b[29]), .c(c[28]));
fa_dataflow g30 (.s(s[30]), .cout(c[30]), .a(a[30]), .b(b[30]), .c(c[29]));
fa_dataflow g31 (.s(s[31]), .cout(cout), .a(a[31]), .b(b[31]), .c(c[30]));

endmodule
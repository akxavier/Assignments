module nor_gate
(output out,
input a, b);

nor g1 (out, a, b);

endmodule 
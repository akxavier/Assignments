module array_of_16_or_gate
(output [15:0] out,
input [15:0] a, b);

or g[15:0] (out, a, b);

endmodule 
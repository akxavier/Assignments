module nand_gate
(output out,
input a, b);

nand g1 (out, a, b);

endmodule
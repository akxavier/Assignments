module or_gate
(output out,
input a, b);

or g1 (out, a, b);

endmodule 